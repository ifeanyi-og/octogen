// src/rtl/octogen_top.v
module octogen_top (
    input  wire clk,
    input  wire rst_n
    // TODO: add ADC / Ethernet / debug I/O later
);


endmodule